module Decodificador #(
    parameter W = 4
) (
    input [W-1:0] i_Display,
    output reg [6:0] o_Display
);

  always @(*) begin
    case (i_Display)
      4'b0000: o_Display <= 7'b1000000;  //0
      4'b0001: o_Display <= 7'b1111001;  //1
      4'b0010: o_Display <= 7'b0100100;  //2
      4'b0011: o_Display <= 7'b0110000;  //3
      4'b0100: o_Display <= 7'b0011001;  //4
      4'b0101: o_Display <= 7'b0010010;  //5
      4'b0110: o_Display <= 7'b0000010;  //6
      4'b0111: o_Display <= 7'b1111000;  //7
      4'b1000: o_Display <= 7'b0000000;  //8
      4'b1001: o_Display <= 7'b0011000;  //9
      4'b1010: o_Display <= 7'b0001000;  //A
      4'b1011: o_Display <= 7'b0000011;  //B
      4'b1100: o_Display <= 7'b1000110;  //C
      4'b1101: o_Display <= 7'b0100001;  //D
      4'b1110: o_Display <= 7'b0000110;  //E
      4'b1111: o_Display <= 7'b0001110;  //F
      default: o_Display <= 7'b1111111;  //resto
    endcase
  end

endmodule